module mruby

#flag -L @VMODROOT/lib
#flag -I @VMODROOT/include/mruby-3.1.0
#flag @VMODROOT/lib/mruby-3.1.0/libmruby.a -lm
