module main

import src.mruby

fn main() {
}
